package my_pkg;
	import uvm_pkg::*;

	`include "my_sequence.sv"
    `include "my_sequencer.sv"
	`include "my_monitor.sv"
	`include "my_driver.sv"
	`include "my_agent.sv"
	`include "my_scoreboard.sv"
    `include "my_config.sv"
	`include "my_env.sv"
	`include "test_pkg.sv"
endpackage