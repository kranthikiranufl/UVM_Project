 package my_pkg;
  import uvm_pkg::*;

 `include "my_sequencer.sv"
 `include "my_driver.sv"
 `include "my_monitor.sv"
 `include "my_agent.sv"
 `include "my_sb.sv"
 `include "my_env.sv"
 `include "my_test.sv"
endpackage
