interface dut_if (input clk);
 logic [7:0] a,b;
 logic  [15:0] c;
endinterface
